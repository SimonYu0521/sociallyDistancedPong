`default_nettype none

// juse SW 17-15 to set the color
// 
// KEY 1 loads the color into the pixel
// KEY 2 displays the colors
module ChipInterface(input logic CLOCK_50, 
		     input logic [3:0] KEY,
		     input logic [17:0] SW,
		     output logic NEO_OUT,
		     output logic [17:0] LEDR);

	logic add_red, add_green, add_blue, reset, load, go, ready; 
	logic [4:0] pixel;
	

	Synchronizer SyncR (.asynchronous(SW[17]), .local_clock(CLOCK_50), .synchronized(add_red));
	Synchronizer SyncG (.asynchronous(SW[16]), .local_clock(CLOCK_50), .synchronized(add_green));
	Synchronizer SyncB (.asynchronous(SW[15]), .local_clock(CLOCK_50), .synchronized(add_blue));
	
	Synchronizer SyncP0 (.asynchronous(SW[0]), .local_clock(CLOCK_50), .synchronized(pixel[0]));
	Synchronizer SyncP1 (.asynchronous(SW[1]), .local_clock(CLOCK_50), .synchronized(pixel[1]));
	Synchronizer SyncP2 (.asynchronous(SW[2]), .local_clock(CLOCK_50), .synchronized(pixel[2]));
   Synchronizer SyncP3 (.asynchronous(SW[3]), .local_clock(CLOCK_50), .synchronized(pixel[3]));
	Synchronizer SyncP4 (.asynchronous(SW[4]), .local_clock(CLOCK_50), .synchronized(pixel[4]));


	Synchronizer SyncK0 (.asynchronous(~KEY[0]), .local_clock(CLOCK_50), .synchronized(reset));
	Synchronizer SyncK1 (.asynchronous(~KEY[1]), .local_clock(CLOCK_50), .synchronized(load));
	Synchronizer SyncK2 (.asynchronous(~KEY[2]), .local_clock(CLOCK_50), .synchronized(go));
	
	

	SetNeopix SN (.neopixel_data(NEO_OUT), .*);
	
	assign LEDR[0] = ready;

endmodule: ChipInterface

	
	

module SetNeopix (input logic add_red, add_green, add_blue, reset, CLOCK_50, 
		  input logic [4:0] pixel,
	    input logic load, go,
		  output logic neopixel_data, ready);

	logic [7:0] red, blue, green;
  logic go_npx;

	NeopixelController NC (.go(go_npx), .*);
  NPX_GO_fsm Ctrl_FSM (.clock(CLOCK_50), .reset_n(~reset), .go, .ready, .go_npx);
	
	assign red = add_red ? 8'hFF : 8'd0;
	assign green = add_green ? 8'hFF : 8'd0;
	assign blue = add_blue ? 8'hff : 8'd0;

  // assign red = add_red ? {3'b0, pixel} : 8'd0;
	// assign green = add_green ? {3'b0, pixel} : 8'd0;
	// assign blue = add_blue ? {3'b0, pixel} : 8'd0;


endmodule: SetNeopix

// Automatically generated by ferris highroller on 2/9/2022, 2:50:28 PM
module NPX_GO_fsm (
  input logic clock, reset_n,
  input logic go,
  input logic ready,
  output logic go_npx
  );
  
  enum logic [1:0] {
    WAIT_GO_AND_READY,
    WAIT_GO_UNASSERT,
    SEND_GO
  } cstate, nstate;
  
  always_comb begin
    nstate = cstate;
    go_npx = 1'b0;
    
    case (cstate)
      WAIT_GO_AND_READY: begin
        if (go & ready) begin
		  go_npx = 1'b1;
          nstate = SEND_GO;
         
        end
      end
      WAIT_GO_UNASSERT: begin
        if (~go) begin
          nstate = WAIT_GO_AND_READY;
        end
      end
      SEND_GO: begin
		 nstate = WAIT_GO_UNASSERT;
        go_npx = 1'b1;
        
      end
    endcase
  end
  always_ff @(posedge clock, negedge reset_n) begin
    if (!reset_n) cstate <= WAIT_GO_AND_READY;
    else cstate <= nstate;
  end
  
endmodule : NPX_GO_fsm